//Basic NOT 
module not (in, out);
input in;
output out;
assign out = ~in;
endmodule

